// This file is part of Small Practice CPU.
// 
// Copyright 2016 by Andrew Clark (FL4SHK).
// 
// Small Practice CPU is free software: you can redistribute it and/or
// modify it under the terms of the GNU General Public License as published
// by the Free Software Foundation, either version 3 of the License, or (at
// your option) any later version.
// 
// Small Practice CPU is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
// 
// You should have received a copy of the GNU General Public License along
// with Small Practice CPU.  If not, see <http://www.gnu.org/licenses/>.


`include "src/alu_defines.svinc"

`include "src/instr_decoder_defines.svinc"
//`include "src/cpu_extras_defines.svinc"


module spcpu_test_bench;
	
	bit clk_gen_reset, tb_clk;
	
	bit test_mem_reset;
	
	//// Various test bench reset signals
	//bit alu_tb_reset, 
	//	instr_grp_dec_tb_reset,
	//	instr_dec_tb_reset;
	
	// reset signal for test_cpu
	bit test_cpu_reset;
	
	
	tb_clk_gen clk_gen( .reset(clk_gen_reset), .clk(tb_clk) );
	
	
	//alu_test_bench alu_tb( .tb_clk(tb_clk), .reset(alu_tb_reset) );
	//instr_group_decoder_test_bench instr_grp_dec_tb( .tb_clk(tb_clk), 
	//	.reset(instr_grp_dec_tb_reset) );
	//instr_decoder_test_bench instr_dec_tb( .tb_clk(tb_clk),
	//	.reset(instr_dec_tb_reset) );
	
	tb_mem_inputs mem_inputs;
	//logic [`cpu_data_inout_16_msb_pos:0] tb_mem_read_data_out ;
	wire [`cpu_data_inout_16_msb_pos:0] tb_mem_read_data_out ;
	
	tb_memory test_mem( .write_clk(tb_clk), .reset(test_mem_reset),
		.the_inputs(mem_inputs), .read_data_out(tb_mem_read_data_out) );
	
	`include "src/test_mem_tasks.svinc"
	
	
	wire [`cpu_data_inout_16_msb_pos:0] test_cpu_data_inout_direct;
	bit [`cpu_addr_msb_pos:0] test_cpu_data_inout_addr;
	bit test_cpu_data_acc_sz, test_cpu_data_inout_we;
	
	spcpu test_cpu( .clk(tb_clk), .reset(test_cpu_reset),
		.data_inout(test_cpu_data_inout_direct),
		.data_inout_addr(test_cpu_data_inout_addr),
		.data_acc_sz(test_cpu_data_acc_sz),
		.data_inout_we(test_cpu_data_inout_we) );
	
	//logic [`cpu_data_inout_16_msb_pos:0] test_cpu_data_in, 
	//	test_cpu_data_out;
	logic [`cpu_data_inout_16_msb_pos:0] test_cpu_data_out;
	
	
	//assign test_cpu_data_inout_direct = (!test_cpu_data_inout_we) 
	//	? test_cpu_data_in : `cpu_data_inout_16_width'hz;
	assign test_cpu_data_inout_direct = (!test_cpu_data_inout_we) 
		? tb_mem_read_data_out : `cpu_data_inout_16_width'hz;
	
	assign test_cpu_data_out = (test_cpu_data_inout_we)
		? test_cpu_data_inout_direct : `cpu_data_inout_16_width'hz;
	
	
	initial
	begin
		clk_gen_reset = 1'b0;
		test_cpu_reset = 1'b0;
		
		{ mem_inputs.write_addr_in, mem_inputs.write_data_in,
			mem_inputs.write_data_acc_sz, mem_inputs.write_data_we } = 0;
		
		#2
		clk_gen_reset = 1'b1;
		test_cpu_reset = 1'b1;
		
		#2
		test_cpu_reset = 1'b0;
		
	end
	
	
	always @ ( posedge tb_clk )
	begin
		
		// If the CPU wants to read or write 8-bit data
		if ( test_cpu_data_acc_sz == pkg_cpu::cpu_data_acc_sz_8 )
		begin
			// If the CPU wants to read 8-bit data
			if (!test_cpu_data_inout_we)
			begin
				read_test_mem_8(test_cpu_data_inout_addr);
				
				//$display( "%h", test_cpu_data_in );
			end
			
			// If the CPU wants to write 8-bit data
			else // if (test_cpu_data_inout_we)
			begin
				write_test_mem_8( test_cpu_data_inout_addr, 
					test_cpu_data_out );
			end
		end
		
		
		// If the CPU wants to read or write 16-bit data
		else // if ( test_cpu_data_acc_sz == pkg_cpu::cpu_data_acc_sz_16 )
		begin
			// If the CPU wants to read 16-bit data (for Small Practice
			// CPU, it's used for loading either a 16-bit instruction or
			// a 16-bit half of a 32-bit instruction)
			if (!test_cpu_data_inout_we)
			begin
				read_test_mem_16(test_cpu_data_inout_addr);
			end
			
			// If the CPU wants to write 16-bit data (which should NOT 
			// happen with the current design of Small Practice CPU)
			else // if (test_cpu_data_inout_we)
			begin
				$display( "spcpu_test_bench:  Uh oh!  The CPU module ",
					"wants to store a 16-bit value!  That should NOT ",
					"happen!" );
			end
		end
		
	end
	
	
endmodule



`define make_reg_pair( index_hi ) `make_pair( cpu_regs, index_hi )

// Make reg pair with pair index
`define make_reg_pair_w_pi( pair_index ) `make_pair( cpu_regs, \
	pair_index << 1 )

`define get_cpu_rp_pc `make_reg_pair_w_pi(pkg_cpu::cpu_rp_pc_pind)
`define get_cpu_rp_lr `make_reg_pair_w_pi(pkg_cpu::cpu_rp_lr_pind)

// The next value of the PC after a non-PC-changing 16-bit instruction, or
// the next value of data_inout_addr after loading the high 16 bits of a
// 32-bit instruction
`define get_pc_after_reg_instr_16 ( `get_cpu_rp_pc + 2 )

// The next value of the PC after a non-PC-changing 32-bit instruction
`define get_pc_after_reg_instr_32 ( `get_cpu_rp_pc + 4 )


`define wire_rhs_pc_indices_contain_reg_index( reg_index ) \
	( ( reg_index == pkg_cpu::cpu_rp_pc_hi_rind ) \
	|| ( reg_index == pkg_cpu::cpu_rp_pc_lo_rind ) )

`define wire_rhs_rp_index_is_pc_index( rp_index ) \
	( rp_index == pkg_cpu:: cpu_rp_pc_pind )


// The CPU itself
module spcpu
	
	import pkg_cpu::*;
	import pkg_pflags::*;
	import pkg_instr_dec::*;
	import pkg_alu::*;
	
	( input bit clk, input bit reset,
	
	// Data being read in or written out
	inout [`cpu_data_inout_16_msb_pos:0] data_inout,
	
	// The address being loaded from or written to
	output bit [`cpu_addr_msb_pos:0] data_inout_addr,
	
	// Size (8-bit or 16-bit) of data being read/written
	output bit data_acc_sz,
	
	// Write enable, which when low specifies that the CPU wants to read,
	// and when high specifies that the CPU wants to write,
	output bit data_inout_we );
	
	
	
	
	
	
	
	// CPU state stuff
	// For some reason, vvp does weird things when I make cpu_regs part of
	// the misc_cpu_vars struct, so just get rid of that struct for now.
	bit [`cpu_reg_msb_pos:0] cpu_regs[0:`cpu_reg_arr_msb_pos];
	
	// The entirety of a 16-bit insturction, or the high 16 bits of a
	// 32-bit instruction
	bit [`instr_main_msb_pos:0] instr_in_hi,
	
	// The low 16 bits of a 32-bit instruction
		instr_in_lo;
	
	// The current CPU state
	bit [`cpu_state_msb_pos:0] curr_state;
	
	// Whether or not the instruction changed the pc
	bit instr_changes_pc;
	
	// These are used for communication with the outside world
	wire [`cpu_data_inout_16_msb_pos:0] temp_data_in;
	bit [`cpu_data_inout_16_msb_pos:0] temp_data_out;
	
	
	`include "src/extra_wires.svinc"
	
	
	
	
	// Instruction decoding struct and enum instances
	
	// The instr_group that is the output of the instr_group_decoder module
	// called instr_grp_dec
	instr_group init_instr_grp;
	
	// The instr_group instance that is used after loading the first 16
	// bits of an instruction
	instr_group final_instr_grp;
	
	ig1_dec_outputs ig1d_outputs;
	ig2_dec_outputs ig2d_outputs;
	ig3_dec_outputs ig3d_outputs;
	ig4_dec_outputs ig4d_outputs;
	ig5_dec_outputs ig5d_outputs;
	
	
	
	// Instruction decoder modules
	instr_group_decoder instr_grp_dec( .instr_hi(temp_data_in),
		.group_out(init_instr_grp) );
	
	instr_grp_1_decoder instr_grp_1_dec( .instr_hi(temp_data_in),
		.ig1d_outputs(ig1d_outputs) );
	instr_grp_2_decoder instr_grp_2_dec( .instr_hi(temp_data_in),
		.ig2d_outputs(ig2d_outputs) );
	instr_grp_3_decoder instr_grp_3_dec( .instr_hi(temp_data_in),
		.ig3d_outputs(ig3d_outputs) );
	instr_grp_4_decoder instr_grp_4_dec( .instr_hi(temp_data_in),
		.ig4d_outputs(ig4d_outputs) );
	instr_grp_5_decoder instr_grp_5_dec( .instr_hi(temp_data_in),
		.ig5d_outputs(ig5d_outputs) );
	
	
	// Outside world access assign statements
	assign data_inout = (data_inout_we) ? temp_data_out
		: `cpu_data_inout_16_width'hz;
	assign temp_data_in = (!data_inout_we) ? data_inout
		: `cpu_data_inout_16_width'hz;
	
	
	
	`include "src/extra_wire_assignments.svinc"
	
	
	
	// Tasks
	`include "src/debug_tasks.svinc"
	
	`include "src/state_changing_tasks.svinc"
	
	`include "src/instr_exec_tasks.svinc"
	
	`include "src/check_instr_changes_pc_tasks.svinc"
	
	
	bit ready;
	initial ready = 0;
	
	always @ ( posedge clk )
	begin
	
	if (reset)
	begin
		//{ data_inout_addr, data_inout_we } = 0;
		data_inout_addr <= 0;
		data_inout_we <= 0;
		
		data_acc_sz <= pkg_cpu::cpu_data_acc_sz_16;
		
		
		// Clear every CPU register
		{ cpu_regs[0], cpu_regs[1], cpu_regs[2], cpu_regs[3], 
			cpu_regs[4], cpu_regs[5], cpu_regs[6], cpu_regs[7],
			cpu_regs[8], cpu_regs[9], cpu_regs[10], cpu_regs[11],
			cpu_regs[12], cpu_regs[13], cpu_regs[14], cpu_regs[15] } <= 0;
		
		curr_state <= pkg_cpu::cpu_st_load_instr_hi;
		
		ready <= 0;
	end
	
	end
	
	
	
	always @ ( posedge clk )
	begin
		if ( `get_cpu_rp_pc >= 20 * 2 )
		begin
			$display("\ndone");
			$finish;
		end
	end
	
	
	
	always @ ( posedge clk )
	begin
		
		//$display( "%h", `get_cpu_rp_pc );
		//$display( "%h", curr_state == pkg_cpu::cpu_st_load_instr_hi );
		
		if (!ready)
		begin
			ready <= 1;
			advance_pc_etc_after_reg_instr_16();
			prepare_to_load_16_no_addr();
		end
		
		else if ( curr_state == pkg_cpu::cpu_st_load_instr_hi )
		begin
			// Back up temp_data_in and init_instr_grp
			instr_in_hi <= temp_data_in;
			final_instr_grp <= init_instr_grp;
			
			if ( init_instr_grp != pkg_instr_dec::instr_grp_5 )
			begin
				//instr_in_hi <= temp_data_in;
				curr_state <= pkg_cpu::cpu_st_start_exec_instr;
			end
			
			// Handle 32-bit instructions
			else if ( init_instr_grp == pkg_instr_dec::instr_grp_5 )
			begin
				//instr_in_hi <= temp_data_in;
				curr_state <= pkg_cpu::cpu_st_load_instr_lo;
				
				advance_dio_addr_for_instr_lo();
				prepare_to_load_16_no_addr();
			end
			
			else // if ( init_instr_grp 
				// == pkg_instr_dec::instr_grp_unknown )
			begin
				$display("Unknown instruction encoding");
				
				//curr_state <= pkg_cpu::cpu_st_load_instr_hi;
			end
			
		end
		
		else if ( curr_state == pkg_cpu::cpu_st_load_instr_lo )
		begin
			curr_state <= pkg_cpu::cpu_st_start_exec_instr;
			instr_in_lo <= temp_data_in;
		end
		
		
		// Instruction execution states
		else if ( curr_state == pkg_cpu::cpu_st_start_exec_instr )
		begin
			start_exec_instr();
		end
		
		else // if ( curr_state == pkg_cpu::cpu_st_finish_exec_instr )
		begin
			finish_exec_instr();
			
			//curr_state <= pkg_cpu::cpu_st_load_instr_hi;
		end
		
	end
	
	
	
	always @ ( curr_state )
	begin
		if ( ready && curr_state == pkg_cpu::cpu_st_load_instr_hi )
		begin
			if ( init_instr_grp == pkg_instr_dec::instr_grp_1 )
			begin
				check_grp_1_instr_for_pc_change();
			end
			
			else if ( init_instr_grp == pkg_instr_dec::instr_grp_2 )
			begin
				check_grp_2_instr_for_pc_change();
			end
			
			else if ( init_instr_grp == pkg_instr_dec::instr_grp_3 )
			begin
				check_grp_3_instr_for_pc_change();
			end
			
			else if ( init_instr_grp == pkg_instr_dec::instr_grp_4 )
			begin
				check_grp_4_instr_for_pc_change();
			end
			
			else if ( init_instr_grp == pkg_instr_dec::instr_grp_5 )
			begin
				check_grp_5_instr_for_pc_change();
			end
			
		end
		
	end
	
	
	
endmodule


