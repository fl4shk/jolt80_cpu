// This file is part of Small Practice CPU.
// 
// Copyright 2016 by Andrew Clark (FL4SHK).
// 
// Small Practice CPU is free software: you can redistribute it and/or
// modify it under the terms of the GNU General Public License as published
// by the Free Software Foundation, either version 3 of the License, or (at
// your option) any later version.
// 
// Small Practice CPU is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
// 
// You should have received a copy of the GNU General Public License along
// with Small Practice CPU.  If not, see <http://www.gnu.org/licenses/>.


`include "src/alu_defines.svinc"

`include "src/instr_decoder_defines.svinc"
//`include "src/cpu_extras_defines.svinc"


module spcpu_test_bench;
	
	bit clk_gen_reset, tb_half_clk, tb_mem_clk;
	
	bit test_mem_reset;
	
	
	// reset signal for test_cpu
	bit test_cpu_reset;
	
	
	tb_half_clk_gen half_clk_gen( .reset(clk_gen_reset), 
		.half_clk(tb_half_clk) );
	tb_memory_clk_gen mem_clk_gen( .reset(clk_gen_reset), 
		.mem_clk(tb_mem_clk) );
	
	
	
	wire [`cpu_data_inout_16_msb_pos:0] tb_mem_read_data_out;
	
	wire [`cpu_data_inout_16_msb_pos:0] test_cpu_data_inout_direct;
	bit [`cpu_addr_msb_pos:0] test_cpu_data_inout_addr;
	bit test_cpu_data_acc_sz, test_cpu_data_inout_we;
	logic [`cpu_data_inout_16_msb_pos:0] test_cpu_data_out;
	
	spcpu test_cpu( .clk(tb_half_clk), .reset(test_cpu_reset),
		.data_inout(test_cpu_data_inout_direct),
		.data_inout_addr(test_cpu_data_inout_addr),
		.data_acc_sz(test_cpu_data_acc_sz),
		.data_inout_we(test_cpu_data_inout_we) );
	
	//tb_memory test_mem( .clk(tb_mem_clk), .reset(test_mem_reset),
	//	.the_inputs(mem_inputs), .read_data_out(tb_mem_read_data_out) );
	tb_memory test_mem( .clk(tb_mem_clk), .reset(test_mem_reset),
		.addr_in(test_cpu_data_inout_addr),
		.write_data_in(test_cpu_data_out),
		.data_acc_sz(test_cpu_data_acc_sz),
		.write_data_we(test_cpu_data_inout_we), 
		.read_data_out(tb_mem_read_data_out) );
	
	
	
	
	
	//assign test_cpu_data_inout_direct = (!test_cpu_data_inout_we) 
	//	? test_cpu_data_in : `cpu_data_inout_16_width'hz;
	assign test_cpu_data_inout_direct = (!test_cpu_data_inout_we) 
		? tb_mem_read_data_out : `cpu_data_inout_16_width'hz;
	//assign test_cpu_data_inout_direct = (!test_cpu_data_inout_we) 
	//	? temp_read_data_out : `cpu_data_inout_16_width'hz;
	
	assign test_cpu_data_out = (test_cpu_data_inout_we)
		? test_cpu_data_inout_direct : `cpu_data_inout_16_width'hz;
	
	
	
	initial
	begin
		clk_gen_reset = 1'b1;
		test_cpu_reset = 1'b0;
		//$display(test_cpu_reset);
		
		#4
		test_cpu_reset = 1'b1;
		//$display(test_cpu_reset);
		
		//{ mem_inputs.write_addr_in, mem_inputs.write_data_in,
		//	mem_inputs.write_data_acc_sz, mem_inputs.write_data_we } = 0;
		
		#4
		test_cpu_reset = 1'b0;
		
	end
	
	//always @ ( posedge tb_half_clk )
	//begin
	//	$display( "%h %h %h %h", test_cpu_data_inout_direct,
	//		test_cpu_data_inout_addr, test_cpu_data_acc_sz, 
	//		test_cpu_data_inout_we );
	//end
	
	
endmodule



`define make_reg_pair( index_hi ) `make_pair( cpu_regs, index_hi )

// Make reg pair with pair index
`define make_reg_pair_w_pi( pair_index ) \
	`make_reg_pair( `make_reg_ind_from_pi(pair_index) )

`define get_cpu_rp_pc `make_reg_pair_w_pi(pkg_cpu::cpu_rp_pc_pind)
`define get_cpu_rp_lr `make_reg_pair_w_pi(pkg_cpu::cpu_rp_lr_pind)



`define instr_16_num_bytes 2
`define instr_32_num_bytes 4

// The next value of the PC after a non-PC-changing 16-bit instruction, or
// the next value of data_inout_addr after loading the high 16 bits of a
// 32-bit instruction
//`define get_pc_after_reg_instr_16 ( `get_cpu_rp_pc + `instr_16_num_bytes )
`define get_pc_after_reg_instr ( `get_cpu_rp_pc + `instr_16_num_bytes )

// The next value of the PC after a non-PC-changing 32-bit instruction
//`define get_pc_after_reg_instr_32 ( `get_cpu_rp_pc + `instr_32_num_bytes )


`define wire_rhs_pc_indices_contain_reg_index( reg_index ) \
	( ( reg_index == pkg_cpu::cpu_rp_pc_hi_rind ) \
	|| ( reg_index == pkg_cpu::cpu_rp_pc_lo_rind ) )
`define wire_rhs_rp_index_is_pc_index( rp_index ) \
	( rp_index == pkg_cpu::cpu_rp_pc_pind )


// The CPU itself
module spcpu
	
	import pkg_cpu::*;
	import pkg_pflags::*;
	import pkg_instr_dec::*;
	import pkg_alu::*;
	
	( input bit clk, input bit reset,
	
	// Data being read in or written out
	inout [`cpu_data_inout_16_msb_pos:0] data_inout,
	
	// The address being loaded from or written to
	output bit [`cpu_addr_msb_pos:0] data_inout_addr,
	
	// Size (8-bit or 16-bit) of data being read/written
	output bit data_acc_sz,
	
	// Write enable, which when low specifies that the CPU wants to read,
	// and when high specifies that the CPU wants to write,
	output bit data_inout_we );
	
	
	
	
	
	
	
	// CPU state stuff
	// For some reason, vvp does weird things when I make cpu_regs part of
	// the misc_cpu_vars struct, so just get rid of that struct for now.
	bit [`cpu_reg_msb_pos:0] cpu_regs[0:`cpu_reg_arr_msb_pos];
	
	bit [ `cpu_reg_width + `cpu_reg_msb_pos : 0 ] prev_pc;
	wire [`cpu_reg_msb_pos:0] prev_r14, prev_r15;
	assign { prev_r14, prev_r15 } = prev_pc;
	
	
	// The entirety of a 16-bit insturction, or the high 16 bits of a
	// 32-bit instruction
	bit [`instr_main_msb_pos:0] instr_in_hi,
	
	// The low 16 bits of a 32-bit instruction
		instr_in_lo;
	
	// The current CPU state
	bit [`cpu_state_msb_pos:0] curr_state;
	
	
	
	// These are used for communication with the outside world
	wire [`cpu_data_inout_16_msb_pos:0] temp_data_in;
	bit [`cpu_data_inout_16_msb_pos:0] temp_data_out;
	
	
	
	
	
	`include "src/extra_instr_dec_vars.svinc"
	`include "src/alu_vars.svinc"
	
	
	
	
	// Instruction decoding struct and enum instances
	
	// The instr_group that is the output of the instr_group_decoder module
	// called instr_grp_dec
	instr_group init_instr_grp;
	
	// The instr_group instance that is used after loading the first 16
	// bits of an instruction
	instr_group final_instr_grp;
	
	
	
	
	// Module instances
	instr_group_decoder instr_grp_dec( .instr_hi(temp_data_in),
		.group_out(init_instr_grp) );
	
	instr_grp_1_decoder instr_grp_1_dec( .instr_hi(temp_data_in),
		.opcode(ig1_opcode), .ra_index(ig1_ra_index),
		.imm_value_8(ig1_imm_value_8),
		.ra_index_is_for_pair(ig1_ra_index_is_for_pair) );
	instr_grp_2_decoder instr_grp_2_dec( .instr_hi(temp_data_in),
		.opcode(ig2_opcode), 
		.ra_index(ig2_ra_index),
		.rb_index(ig2_rb_index),
		.ra_index_is_for_pair(ig2_ra_index_is_for_pair),
		.rb_index_is_for_pair(ig2_rb_index_is_for_pair) );
	instr_grp_3_decoder instr_grp_3_dec( .instr_hi(temp_data_in),
		.opcode(ig3_opcode), 
		.ra_index(ig3_ra_index),
		.rbp_index(ig3_rbp_index), 
		.rcp_index(ig3_rcp_index) );
	instr_grp_4_decoder instr_grp_4_dec( .instr_hi(temp_data_in),
		.opcode(ig4_opcode), 
		.imm_value_8(ig4_imm_value_8) );
	instr_grp_5_decoder instr_grp_5_dec( .instr_hi(temp_data_in),
		.opcode(ig5_opcode), 
		.ra_index(ig5_ra_index),
		.rbp_index(ig5_rbp_index),
		.ra_index_is_for_pair(ig5_ra_index_is_for_pair) );
	
	alu the_alu( .oper(the_alu_op), .a_in_hi(alu_a_in_hi),
		.a_in_lo(alu_a_in_lo), .b_in(alu_b_in), 
		.proc_flags_in(alu_proc_flags_in), .out_hi(alu_out_hi),
		.out_lo(alu_out_lo), .proc_flags_out(alu_proc_flags_out) );
	
	
	// Outside world access assign statements
	assign data_inout = (data_inout_we) ? temp_data_out
		: `cpu_data_inout_16_width'hz;
	assign temp_data_in = (!data_inout_we) ? data_inout
		: `cpu_data_inout_16_width'hz;
	
	
	
	
	
	
	`include "src/extra_wire_assignments.svinc"
	
	
	
	// Tasks
	`include "src/debug_tasks.svinc"
	
	`include "src/state_changing_tasks.svinc"
	
	`include "src/update_instr_possibly_changes_pc_tasks.svinc"
	
	`include "src/extra_instr_dec_tasks_funcs.svinc"
	
	`include "src/debug_disassembly_tasks.svinc"
	
	`include "src/instr_exec_tasks.svinc"
	
	`include "src/alu_control_tasks.svinc"
	
	
	bit ready;
	initial ready = 0;
	
	
	// This is used to determine when to stop simulation
	logic [5:0] data_in_is_0_counter;
	
	always @ ( posedge clk )
	begin
	
	if (reset)
	begin
		//{ data_inout_addr, data_inout_we } <= 0;
		data_inout_addr <= 0;
		data_inout_we <= 0;
		
		data_acc_sz <= pkg_cpu::cpu_data_acc_sz_16;
		
		
		// Clear every CPU register
		{ cpu_regs[0], cpu_regs[1], cpu_regs[2], cpu_regs[3], 
			cpu_regs[4], cpu_regs[5], cpu_regs[6], cpu_regs[7],
			cpu_regs[8], cpu_regs[9], cpu_regs[10], cpu_regs[11],
			cpu_regs[12], cpu_regs[13], cpu_regs[14], cpu_regs[15] } <= 0;
		
		//curr_state <= pkg_cpu::cpu_st_begin_0;
		curr_state <= 0;
		ready <= 1;
		
		data_in_is_0_counter <= 0;
		
		prep_load_16_no_addr();
	end
	
	end
	
	
	
	// End CPU simulation if there are a bunch of 0000's in a row
	always @ ( posedge clk )
	begin
		if ( curr_state == pkg_cpu::cpu_st_load_instr_hi )
		begin
			if ( temp_data_in == 0 )
			begin
				data_in_is_0_counter <= data_in_is_0_counter + 1;
			end
			
			else
			begin
				data_in_is_0_counter <= 0;
			end
			
			if ( data_in_is_0_counter >= 4 )
			begin
				$display("\ndone");
				$finish;
			end
		end
	end
	
	
	always @ ( posedge clk )
	begin
	
	if (ready)
	begin
		if ( curr_state == pkg_cpu::cpu_st_begin_0 )
		begin
			curr_state <= curr_state + 1;
			prep_load_16_no_addr();
		end
		
		
		else if ( curr_state == pkg_cpu::cpu_st_load_instr_hi )
		begin
			debug_disp_regs_and_proc_flags();
			$display();
			
			
			// Back up temp_data_in, init_instr_grp, and pc
			instr_in_hi <= temp_data_in;
			final_instr_grp <= init_instr_grp;
			prev_pc <= `get_cpu_rp_pc;
			
			
			// Back up the decoded instruction contents to be used on
			// cycles after the current one.
			back_up_ig1_instr_contents();
			back_up_ig2_instr_contents();
			back_up_ig3_instr_contents();
			back_up_ig4_instr_contents();
			back_up_ig5_instr_contents();
			
			update_extra_ig1_pc_stuff();
			update_extra_ig2_pc_stuff();
			update_extra_ig3_pc_stuff();
			//update_extra_ig4_pc_stuff();
			update_extra_ig5_pc_stuff();
			
			
			
			//if ( init_instr_grp != pkg_instr_dec::instr_grp_5 )
			if (!init_instr_is_32_bit)
			begin
				curr_state <= pkg_cpu::cpu_st_start_exec_instr;
				
				prep_alu_if_needed_init();
				
			end
			
			// Handle 32-bit instructions
			else if ( init_instr_grp == pkg_instr_dec::instr_grp_5 )
			begin
				prep_load_instr_lo_reg();
			end
			
			//else if ( init_instr_grp == pkg_instr_dec::instr_grp_... )
			//begin
			//	
			//end
			
			
			else // if ( init_instr_grp 
				// == pkg_instr_dec::instr_grp_unknown )
			begin
				$display("Unknown instruction encoding");
				
			end
			
		end
		
		else if ( curr_state == pkg_cpu::cpu_st_load_instr_lo )
		begin
			curr_state <= pkg_cpu::cpu_st_start_exec_instr;
			instr_in_lo <= temp_data_in;
			prep_alu_if_needed_final();
		end
		
		
		// Instruction execution states
		else if ( curr_state == pkg_cpu::cpu_st_start_exec_instr )
		begin
			start_exec_instr();
		end
		
		else if ( curr_state == pkg_cpu::cpu_st_finish_exec_ldst_instr )
		begin
			finish_exec_ldst_instr();
		end
		
		else // if ( curr_state 
			// == pkg_cpu::cpu_st_update_pc_after_instr_possibly_changed )
		begin
			$display( "Check whether the pc was actually changed by a ",
				 "non-branch, non-call instruction" );
			
			
			// Check if the pc was ACTUALLY changed
			if ( prev_pc == `get_cpu_rp_pc )
			begin
				$display("The pc was not actually changed");
			end
			
			else
			begin
				$display("The pc WAS changed");
			end
			
			prep_load_instr_hi_generic();
			
		end
		
	end
	
	end
	
	
	
	// Combinational logic for updating instr_possibly_changes_pc
	always @ (*)
	begin
		if ( curr_state == pkg_cpu::cpu_st_start_exec_instr )
		begin
			{ instr_is_branch_or_call, non_bc_instr_possibly_changes_pc }
				= 0;
			
			if ( final_instr_grp == pkg_instr_dec::instr_grp_1 )
			begin
				update_ipc_pc_for_grp_1_instr();
			end
			
			else if ( final_instr_grp == pkg_instr_dec::instr_grp_2 )
			begin
				update_ipc_pc_for_grp_2_instr();
			end
			
			else if ( final_instr_grp == pkg_instr_dec::instr_grp_3 )
			begin
				update_ipc_pc_for_grp_3_instr();
			end
			
			else if ( final_instr_grp == pkg_instr_dec::instr_grp_4 )
			begin
				update_ipc_pc_for_grp_4_instr();
			end
			
			else if ( final_instr_grp == pkg_instr_dec::instr_grp_5 )
			begin
				update_ipc_pc_for_grp_5_instr();
			end
		end
	end
	
	
	
endmodule


